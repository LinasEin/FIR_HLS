// ----------------------------------------------------------------------------
// LegUp High-Level Synthesis Tool Version 8.1 (http://www.legupcomputing.com)
// Copyright (c) 2015-2020 LegUp Computing Inc. All Rights Reserved.
// For technical issues, please contact: support@legupcomputing.com
// For general inquiries, please contact: info@legupcomputing.com
// Date: Sat Dec  5 14:04:39 2020
// ----------------------------------------------------------------------------
`define MEMORY_CONTROLLER_ADDR_SIZE 32
// This directory contains the memory initialization files generated by LegUp.
// This relative path is used by ModelSim and FPGA synthesis tool.
`define MEM_INIT_DIR "../mem_init/"

`timescale 1 ns / 1 ns
module FIRFilterStreaming_top
(
	clk,
	reset,
	start,
	finish,
	input_fifo_data_from_source,
	input_fifo_ready_to_source,
	input_fifo_valid_from_source,
	output_fifo_data_to_sink,
	output_fifo_ready_from_sink,
	output_fifo_valid_to_sink
);

input  clk;
input  reset;
input  start;
output reg  finish;
input [31:0] input_fifo_data_from_source;
output reg  input_fifo_ready_to_source;
input  input_fifo_valid_from_source;
output reg [31:0] output_fifo_data_to_sink;
input  output_fifo_ready_from_sink;
output reg  output_fifo_valid_to_sink;
reg  FIRFilterStreaming_inst_clk;
reg  FIRFilterStreaming_inst_reset;
reg  FIRFilterStreaming_inst_start;
wire  FIRFilterStreaming_inst_finish;
reg [31:0] FIRFilterStreaming_inst_input_fifo_data_from_source;
wire  FIRFilterStreaming_inst_input_fifo_ready_to_source;
reg  FIRFilterStreaming_inst_input_fifo_valid_from_source;
wire [31:0] FIRFilterStreaming_inst_output_fifo_data_to_sink;
reg  FIRFilterStreaming_inst_output_fifo_ready_from_sink;
wire  FIRFilterStreaming_inst_output_fifo_valid_to_sink;
reg  FIRFilterStreaming_inst_finish_reg;


FIRFilterStreaming FIRFilterStreaming_inst (
	.clk (FIRFilterStreaming_inst_clk),
	.reset (FIRFilterStreaming_inst_reset),
	.start (FIRFilterStreaming_inst_start),
	.finish (FIRFilterStreaming_inst_finish),
	.input_fifo_data_from_source (FIRFilterStreaming_inst_input_fifo_data_from_source),
	.input_fifo_ready_to_source (FIRFilterStreaming_inst_input_fifo_ready_to_source),
	.input_fifo_valid_from_source (FIRFilterStreaming_inst_input_fifo_valid_from_source),
	.output_fifo_data_to_sink (FIRFilterStreaming_inst_output_fifo_data_to_sink),
	.output_fifo_ready_from_sink (FIRFilterStreaming_inst_output_fifo_ready_from_sink),
	.output_fifo_valid_to_sink (FIRFilterStreaming_inst_output_fifo_valid_to_sink)
);



always @(*) begin
	FIRFilterStreaming_inst_clk = clk;
end
always @(*) begin
	FIRFilterStreaming_inst_reset = reset;
end
always @(*) begin
	FIRFilterStreaming_inst_start = start;
end
always @(*) begin
	FIRFilterStreaming_inst_input_fifo_data_from_source = input_fifo_data_from_source;
end
always @(*) begin
	FIRFilterStreaming_inst_input_fifo_valid_from_source = input_fifo_valid_from_source;
end
always @(*) begin
	FIRFilterStreaming_inst_output_fifo_ready_from_sink = output_fifo_ready_from_sink;
end
always @(posedge clk) begin
	if ((reset | FIRFilterStreaming_inst_start)) begin
		FIRFilterStreaming_inst_finish_reg <= 1'd0;
	end
	if (FIRFilterStreaming_inst_finish) begin
		FIRFilterStreaming_inst_finish_reg <= 1'd1;
	end
end
always @(*) begin
	finish = FIRFilterStreaming_inst_finish;
end
always @(*) begin
	input_fifo_ready_to_source = FIRFilterStreaming_inst_input_fifo_ready_to_source;
end
always @(*) begin
	output_fifo_data_to_sink = FIRFilterStreaming_inst_output_fifo_data_to_sink;
end
always @(*) begin
	output_fifo_valid_to_sink = FIRFilterStreaming_inst_output_fifo_valid_to_sink;
end

endmodule
`timescale 1 ns / 1 ns
module FIRFilterStreaming
(
	clk,
	reset,
	start,
	finish,
	input_fifo_data_from_source,
	input_fifo_ready_to_source,
	input_fifo_valid_from_source,
	output_fifo_data_to_sink,
	output_fifo_ready_from_sink,
	output_fifo_valid_to_sink
);

input  clk;
input  reset;
input  start;
output reg  finish;
input [31:0] input_fifo_data_from_source;
output reg  input_fifo_ready_to_source;
input  input_fifo_valid_from_source;
output reg [31:0] output_fifo_data_to_sink;
input  output_fifo_ready_from_sink;
output reg  output_fifo_valid_to_sink;
reg [31:0] FIRFilterStreaming_entry_0;
reg [31:0] FIRFilterStreaming_entry_1;
reg [31:0] FIRFilterStreaming_entry_2;
reg [30:0] FIRFilterStreaming_entry_bit_select37;
reg [31:0] FIRFilterStreaming_entry_3;
reg [30:0] FIRFilterStreaming_entry_bit_select35;
reg [31:0] FIRFilterStreaming_entry_4;
reg [29:0] FIRFilterStreaming_entry_bit_select33;
reg [31:0] FIRFilterStreaming_entry_5;
reg [29:0] FIRFilterStreaming_entry_bit_select31;
reg [31:0] FIRFilterStreaming_entry_6;
reg [30:0] FIRFilterStreaming_entry_bit_select29;
reg [29:0] FIRFilterStreaming_entry_bit_select27;
reg [31:0] FIRFilterStreaming_entry_7;
reg [28:0] FIRFilterStreaming_entry_bit_select25;
reg [31:0] FIRFilterStreaming_entry_8;
reg [28:0] FIRFilterStreaming_entry_bit_select23;
reg [31:0] FIRFilterStreaming_entry_9;
reg [28:0] FIRFilterStreaming_entry_bit_select21;
reg [31:0] FIRFilterStreaming_entry_10;
reg [30:0] FIRFilterStreaming_entry_bit_select19;
reg [28:0] FIRFilterStreaming_entry_bit_select17;
reg [31:0] FIRFilterStreaming_entry_11;
reg [30:0] FIRFilterStreaming_entry_bit_select15;
reg [28:0] FIRFilterStreaming_entry_bit_select13;
reg [31:0] FIRFilterStreaming_entry_12;
reg [29:0] FIRFilterStreaming_entry_bit_select11;
reg [28:0] FIRFilterStreaming_entry_bit_select9;
reg [31:0] FIRFilterStreaming_entry_13;
reg [29:0] FIRFilterStreaming_entry_bit_select7;
reg [28:0] FIRFilterStreaming_entry_bit_select5;
reg [31:0] FIRFilterStreaming_entry_14;
reg [27:0] FIRFilterStreaming_entry_bit_select1;
reg [31:0] FIRFilterStreaming_entry_15;
reg [27:0] FIRFilterStreaming_entry_bit_select;
reg [31:0] FIRFilterStreaming_entry_bit_concat38;
reg [31:0] FIRFilterStreaming_entry_add_2;
reg [31:0] FIRFilterStreaming_entry_bit_concat36;
reg [31:0] FIRFilterStreaming_entry_sr_add1;
reg [31:0] FIRFilterStreaming_entry_bit_concat34;
reg [31:0] FIRFilterStreaming_entry_newEarly_add_4;
reg [31:0] FIRFilterStreaming_entry_bit_concat32;
reg [31:0] FIRFilterStreaming_entry_sr_add3;
reg [31:0] FIRFilterStreaming_entry_newEarly_add_5;
reg [31:0] FIRFilterStreaming_entry_bit_concat30;
reg [31:0] FIRFilterStreaming_entry_bit_concat28;
reg [31:0] FIRFilterStreaming_entry_sr_add6;
reg [31:0] FIRFilterStreaming_entry_sr_negate;
reg [31:0] FIRFilterStreaming_entry_bit_concat26;
reg [31:0] FIRFilterStreaming_entry_sr_add8;
reg [31:0] FIRFilterStreaming_entry_bit_concat24;
reg [31:0] FIRFilterStreaming_entry_newEarly_newEarly_add_8;
reg [31:0] FIRFilterStreaming_entry_bit_concat22;
reg [31:0] FIRFilterStreaming_entry_sr_add10;
reg [31:0] FIRFilterStreaming_entry_newEarly_newEarly_add_9;
reg [31:0] FIRFilterStreaming_entry_bit_concat20;
reg [31:0] FIRFilterStreaming_entry_bit_concat18;
reg [31:0] FIRFilterStreaming_entry_sr_add13;
reg [31:0] FIRFilterStreaming_entry_bit_concat16;
reg [31:0] FIRFilterStreaming_entry_bit_concat14;
reg [31:0] FIRFilterStreaming_entry_sr_add17;
reg [31:0] FIRFilterStreaming_entry_sr_add18;
reg [31:0] FIRFilterStreaming_entry_bit_concat12;
reg [31:0] FIRFilterStreaming_entry_bit_concat10;
reg [31:0] FIRFilterStreaming_entry_sr_add21;
reg [31:0] FIRFilterStreaming_entry_newEarly_newEarly_add_12;
reg [31:0] FIRFilterStreaming_entry_bit_concat8;
reg [31:0] FIRFilterStreaming_entry_bit_concat6;
reg [31:0] FIRFilterStreaming_entry_sr_add24;
reg [31:0] FIRFilterStreaming_entry_sr_add25;
reg [31:0] FIRFilterStreaming_entry_newEarly_newEarly_add_13;
reg [31:0] FIRFilterStreaming_entry_sr_negate24;
reg [30:0] FIRFilterStreaming_entry_bit_select3;
reg [31:0] FIRFilterStreaming_entry_bit_concat4;
reg [31:0] FIRFilterStreaming_entry_bit_concat2;
reg [31:0] FIRFilterStreaming_entry_sr_add27;
reg [31:0] FIRFilterStreaming_entry_newEarly_newEarly_newEarl;
reg [31:0] FIRFilterStreaming_entry_newCurOp_newEarly_newEarl;
reg [31:0] FIRFilterStreaming_entry_newCurOp_newEarly_add_14;
reg [31:0] FIRFilterStreaming_entry_sr_negate26;
reg [31:0] FIRFilterStreaming_entry_bit_concat;
reg [31:0] FIRFilterStreaming_entry_sr_add28;
reg [31:0] FIRFilterStreaming_entry_newEarly_newEarly_newEarl_var0;
reg [31:0] FIRFilterStreaming_entry_newCurOp_newEarly_newEarl_var1;
reg [31:0] FIRFilterStreaming_entry_newCurOp_newEarly_add_15;
reg [31:0] FIRFilterStreaming_entry_newCurOp_add_15;
reg  FIRFilterStreaming_entry_cmp13;
reg [31:0] FIRFilterStreaming_entry_cond;
reg [31:0] FIRFilterStreaming_previous_0_inferred_reg;
reg [31:0] FIRFilterStreaming_previous_1_inferred_reg;
reg [31:0] FIRFilterStreaming_previous_2_inferred_reg;
reg [31:0] FIRFilterStreaming_previous_3_inferred_reg;
reg [31:0] FIRFilterStreaming_previous_4_inferred_reg;
reg [31:0] FIRFilterStreaming_previous_5_inferred_reg;
reg [31:0] FIRFilterStreaming_previous_6_inferred_reg;
reg [31:0] FIRFilterStreaming_previous_7_inferred_reg;
reg [31:0] FIRFilterStreaming_previous_8_inferred_reg;
reg [31:0] FIRFilterStreaming_previous_9_inferred_reg;
reg [31:0] FIRFilterStreaming_previous_10_inferred_reg;
reg [31:0] FIRFilterStreaming_previous_11_inferred_reg;
reg [31:0] FIRFilterStreaming_previous_12_inferred_reg;
reg [31:0] FIRFilterStreaming_previous_13_inferred_reg;
reg [31:0] FIRFilterStreaming_previous_14_inferred_reg;
reg  FIRFilterStreaming_valid_bit_0;
reg  FIRFilterStreaming_state_stall_0;
reg  FIRFilterStreaming_state_enable_0;
reg  FIRFilterStreaming_valid_bit_1;
reg  FIRFilterStreaming_state_stall_1;
reg  FIRFilterStreaming_state_enable_1;
reg  FIRFilterStreaming_valid_bit_2;
reg  FIRFilterStreaming_state_stall_2;
reg  FIRFilterStreaming_state_enable_2;
reg  FIRFilterStreaming_valid_bit_3;
reg  FIRFilterStreaming_state_stall_3;
reg  FIRFilterStreaming_state_enable_3;
reg  FIRFilterStreaming_II_counter;
reg [31:0] FIRFilterStreaming_entry_newEarly_add_4_reg_stage1;
reg [31:0] FIRFilterStreaming_entry_newEarly_add_5_reg_stage1;
reg [31:0] FIRFilterStreaming_entry_sr_add8_reg_stage1;
reg [31:0] FIRFilterStreaming_entry_newEarly_newEarly_add_8_reg_stage1;
reg [31:0] FIRFilterStreaming_entry_sr_add10_reg_stage1;
reg [31:0] FIRFilterStreaming_entry_sr_add13_reg_stage1;
reg [31:0] FIRFilterStreaming_entry_sr_add18_reg_stage1;
reg [31:0] FIRFilterStreaming_entry_sr_add21_reg_stage1;
reg [31:0] FIRFilterStreaming_entry_newEarly_newEarly_add_12_reg_stage2;
reg [31:0] FIRFilterStreaming_entry_sr_add25_reg_stage1;
reg [31:0] FIRFilterStreaming_entry_newEarly_newEarly_add_13_reg_stage2;
reg [31:0] FIRFilterStreaming_entry_sr_add27_reg_stage1;
reg [31:0] FIRFilterStreaming_entry_newCurOp_newEarly_newEarl_reg_stage2;
reg [31:0] FIRFilterStreaming_entry_sr_add28_reg_stage1;
reg [31:0] FIRFilterStreaming_entry_newCurOp_newEarly_newEarl_var1_reg_stage2;
reg [31:0] FIRFilterStreaming_entry_newCurOp_add_15_reg_stage3;
reg  FIRFilterStreaming_entry_cmp13_reg_stage1;
reg  FIRFilterStreaming_entry_cmp13_reg_stage2;
reg  FIRFilterStreaming_entry_cmp13_reg_stage3;
reg  input_fifo_consumed_valid;
reg [31:0] input_fifo_consumed_data;
reg  input_fifo_consumed_taken;
wire  FIRFilterStreaming_entry_bit_concat38_bit_select_operand_2;
wire  FIRFilterStreaming_entry_bit_concat36_bit_select_operand_2;
wire [1:0] FIRFilterStreaming_entry_bit_concat34_bit_select_operand_2;
wire [1:0] FIRFilterStreaming_entry_bit_concat32_bit_select_operand_2;
wire  FIRFilterStreaming_entry_bit_concat30_bit_select_operand_2;
wire [1:0] FIRFilterStreaming_entry_bit_concat28_bit_select_operand_2;
wire [2:0] FIRFilterStreaming_entry_bit_concat26_bit_select_operand_2;
wire [2:0] FIRFilterStreaming_entry_bit_concat24_bit_select_operand_2;
wire [2:0] FIRFilterStreaming_entry_bit_concat22_bit_select_operand_2;
wire  FIRFilterStreaming_entry_bit_concat20_bit_select_operand_2;
wire [2:0] FIRFilterStreaming_entry_bit_concat18_bit_select_operand_2;
wire  FIRFilterStreaming_entry_bit_concat16_bit_select_operand_2;
wire [2:0] FIRFilterStreaming_entry_bit_concat14_bit_select_operand_2;
wire [1:0] FIRFilterStreaming_entry_bit_concat12_bit_select_operand_2;
wire [2:0] FIRFilterStreaming_entry_bit_concat10_bit_select_operand_2;
wire [1:0] FIRFilterStreaming_entry_bit_concat8_bit_select_operand_2;
wire [2:0] FIRFilterStreaming_entry_bit_concat6_bit_select_operand_2;
wire  FIRFilterStreaming_entry_bit_concat4_bit_select_operand_2;
wire [3:0] FIRFilterStreaming_entry_bit_concat2_bit_select_operand_2;
wire [3:0] FIRFilterStreaming_entry_bit_concat_bit_select_operand_2;
reg  output_fifo_FIRFilterStreaming_state_3_not_accessed_due_to_stall_a;
reg  output_fifo_FIRFilterStreaming_state_3_stalln_reg;
reg  output_fifo_FIRFilterStreaming_state_3_enable_cond_a;


/* Unsynthesizable Statements */
/* synthesis translate_off */
always @(posedge clk)
begin
	if (FIRFilterStreaming_state_enable_0) begin
		$write("FIRFilterStreaming input: %d\n", $signed(FIRFilterStreaming_entry_15));
		// to fix quartus warning
		if (reset == 1'b0 && ^(FIRFilterStreaming_entry_15) === 1'bX) finish <= 0;
	end
	if (FIRFilterStreaming_state_enable_3) begin
		$write("FIRFilterStreaming output: %d\n", $signed(FIRFilterStreaming_entry_cond));
		// to fix quartus warning
		if (reset == 1'b0 && ^(FIRFilterStreaming_entry_cond) === 1'bX) finish <= 0;
	end
end
/* synthesis translate_on */
always @(*) begin
		FIRFilterStreaming_entry_0 = FIRFilterStreaming_previous_14_inferred_reg;
end
always @(*) begin
		FIRFilterStreaming_entry_1 = FIRFilterStreaming_previous_13_inferred_reg;
end
always @(*) begin
		FIRFilterStreaming_entry_2 = FIRFilterStreaming_previous_12_inferred_reg;
end
always @(*) begin
		FIRFilterStreaming_entry_bit_select37 = FIRFilterStreaming_entry_2[30:0];
end
always @(*) begin
		FIRFilterStreaming_entry_3 = FIRFilterStreaming_previous_11_inferred_reg;
end
always @(*) begin
		FIRFilterStreaming_entry_bit_select35 = FIRFilterStreaming_entry_3[30:0];
end
always @(*) begin
		FIRFilterStreaming_entry_4 = FIRFilterStreaming_previous_10_inferred_reg;
end
always @(*) begin
		FIRFilterStreaming_entry_bit_select33 = FIRFilterStreaming_entry_4[29:0];
end
always @(*) begin
		FIRFilterStreaming_entry_5 = FIRFilterStreaming_previous_9_inferred_reg;
end
always @(*) begin
		FIRFilterStreaming_entry_bit_select31 = FIRFilterStreaming_entry_5[29:0];
end
always @(*) begin
		FIRFilterStreaming_entry_6 = FIRFilterStreaming_previous_8_inferred_reg;
end
always @(*) begin
		FIRFilterStreaming_entry_bit_select29 = FIRFilterStreaming_entry_6[30:0];
end
always @(*) begin
		FIRFilterStreaming_entry_bit_select27 = FIRFilterStreaming_entry_6[29:0];
end
always @(*) begin
		FIRFilterStreaming_entry_7 = FIRFilterStreaming_previous_7_inferred_reg;
end
always @(*) begin
		FIRFilterStreaming_entry_bit_select25 = FIRFilterStreaming_entry_7[28:0];
end
always @(*) begin
		FIRFilterStreaming_entry_8 = FIRFilterStreaming_previous_6_inferred_reg;
end
always @(*) begin
		FIRFilterStreaming_entry_bit_select23 = FIRFilterStreaming_entry_8[28:0];
end
always @(*) begin
		FIRFilterStreaming_entry_9 = FIRFilterStreaming_previous_5_inferred_reg;
end
always @(*) begin
		FIRFilterStreaming_entry_bit_select21 = FIRFilterStreaming_entry_9[28:0];
end
always @(*) begin
		FIRFilterStreaming_entry_10 = FIRFilterStreaming_previous_4_inferred_reg;
end
always @(*) begin
		FIRFilterStreaming_entry_bit_select19 = FIRFilterStreaming_entry_10[30:0];
end
always @(*) begin
		FIRFilterStreaming_entry_bit_select17 = FIRFilterStreaming_entry_10[28:0];
end
always @(*) begin
		FIRFilterStreaming_entry_11 = FIRFilterStreaming_previous_3_inferred_reg;
end
always @(*) begin
		FIRFilterStreaming_entry_bit_select15 = FIRFilterStreaming_entry_11[30:0];
end
always @(*) begin
		FIRFilterStreaming_entry_bit_select13 = FIRFilterStreaming_entry_11[28:0];
end
always @(*) begin
		FIRFilterStreaming_entry_12 = FIRFilterStreaming_previous_2_inferred_reg;
end
always @(*) begin
		FIRFilterStreaming_entry_bit_select11 = FIRFilterStreaming_entry_12[29:0];
end
always @(*) begin
		FIRFilterStreaming_entry_bit_select9 = FIRFilterStreaming_entry_12[28:0];
end
always @(*) begin
		FIRFilterStreaming_entry_13 = FIRFilterStreaming_previous_1_inferred_reg;
end
always @(*) begin
		FIRFilterStreaming_entry_bit_select7 = FIRFilterStreaming_entry_13[29:0];
end
always @(*) begin
		FIRFilterStreaming_entry_bit_select5 = FIRFilterStreaming_entry_13[28:0];
end
always @(*) begin
		FIRFilterStreaming_entry_14 = FIRFilterStreaming_previous_0_inferred_reg;
end
always @(*) begin
		FIRFilterStreaming_entry_bit_select1 = FIRFilterStreaming_entry_14[27:0];
end
always @(*) begin
	FIRFilterStreaming_entry_15 = input_fifo_consumed_data;
end
always @(*) begin
		FIRFilterStreaming_entry_bit_select = FIRFilterStreaming_entry_15[27:0];
end
always @(*) begin
		FIRFilterStreaming_entry_bit_concat38 = {FIRFilterStreaming_entry_bit_select37[30:0], FIRFilterStreaming_entry_bit_concat38_bit_select_operand_2};
end
always @(*) begin
		FIRFilterStreaming_entry_add_2 = (FIRFilterStreaming_entry_bit_concat38 + FIRFilterStreaming_entry_1);
end
always @(*) begin
		FIRFilterStreaming_entry_bit_concat36 = {FIRFilterStreaming_entry_bit_select35[30:0], FIRFilterStreaming_entry_bit_concat36_bit_select_operand_2};
end
always @(*) begin
		FIRFilterStreaming_entry_sr_add1 = (FIRFilterStreaming_entry_3 + FIRFilterStreaming_entry_bit_concat36);
end
always @(*) begin
		FIRFilterStreaming_entry_bit_concat34 = {FIRFilterStreaming_entry_bit_select33[29:0], FIRFilterStreaming_entry_bit_concat34_bit_select_operand_2[1:0]};
end
always @(*) begin
		FIRFilterStreaming_entry_newEarly_add_4 = (FIRFilterStreaming_entry_sr_add1 + FIRFilterStreaming_entry_bit_concat34);
end
always @(*) begin
		FIRFilterStreaming_entry_bit_concat32 = {FIRFilterStreaming_entry_bit_select31[29:0], FIRFilterStreaming_entry_bit_concat32_bit_select_operand_2[1:0]};
end
always @(*) begin
		FIRFilterStreaming_entry_sr_add3 = (FIRFilterStreaming_entry_5 + FIRFilterStreaming_entry_bit_concat32);
end
always @(*) begin
		FIRFilterStreaming_entry_newEarly_add_5 = (FIRFilterStreaming_entry_add_2 + FIRFilterStreaming_entry_sr_add3);
end
always @(*) begin
		FIRFilterStreaming_entry_bit_concat30 = {FIRFilterStreaming_entry_bit_select29[30:0], FIRFilterStreaming_entry_bit_concat30_bit_select_operand_2};
end
always @(*) begin
		FIRFilterStreaming_entry_bit_concat28 = {FIRFilterStreaming_entry_bit_select27[29:0], FIRFilterStreaming_entry_bit_concat28_bit_select_operand_2[1:0]};
end
always @(*) begin
		FIRFilterStreaming_entry_sr_add6 = (FIRFilterStreaming_entry_bit_concat30 + FIRFilterStreaming_entry_bit_concat28);
end
always @(*) begin
		FIRFilterStreaming_entry_sr_negate = (32'd0 - FIRFilterStreaming_entry_7);
end
always @(*) begin
		FIRFilterStreaming_entry_bit_concat26 = {FIRFilterStreaming_entry_bit_select25[28:0], FIRFilterStreaming_entry_bit_concat26_bit_select_operand_2[2:0]};
end
always @(*) begin
		FIRFilterStreaming_entry_sr_add8 = (FIRFilterStreaming_entry_sr_negate + FIRFilterStreaming_entry_bit_concat26);
end
always @(*) begin
		FIRFilterStreaming_entry_bit_concat24 = {FIRFilterStreaming_entry_bit_select23[28:0], FIRFilterStreaming_entry_bit_concat24_bit_select_operand_2[2:0]};
end
always @(*) begin
		FIRFilterStreaming_entry_newEarly_newEarly_add_8 = (FIRFilterStreaming_entry_sr_add6 + FIRFilterStreaming_entry_bit_concat24);
end
always @(*) begin
		FIRFilterStreaming_entry_bit_concat22 = {FIRFilterStreaming_entry_bit_select21[28:0], FIRFilterStreaming_entry_bit_concat22_bit_select_operand_2[2:0]};
end
always @(*) begin
		FIRFilterStreaming_entry_sr_add10 = (FIRFilterStreaming_entry_9 + FIRFilterStreaming_entry_bit_concat22);
end
always @(*) begin
		FIRFilterStreaming_entry_newEarly_newEarly_add_9 = (FIRFilterStreaming_entry_sr_add8_reg_stage1 + FIRFilterStreaming_entry_sr_add10_reg_stage1);
end
always @(*) begin
		FIRFilterStreaming_entry_bit_concat20 = {FIRFilterStreaming_entry_bit_select19[30:0], FIRFilterStreaming_entry_bit_concat20_bit_select_operand_2};
end
always @(*) begin
		FIRFilterStreaming_entry_bit_concat18 = {FIRFilterStreaming_entry_bit_select17[28:0], FIRFilterStreaming_entry_bit_concat18_bit_select_operand_2[2:0]};
end
always @(*) begin
		FIRFilterStreaming_entry_sr_add13 = (FIRFilterStreaming_entry_bit_concat20 + FIRFilterStreaming_entry_bit_concat18);
end
always @(*) begin
		FIRFilterStreaming_entry_bit_concat16 = {FIRFilterStreaming_entry_bit_select15[30:0], FIRFilterStreaming_entry_bit_concat16_bit_select_operand_2};
end
always @(*) begin
		FIRFilterStreaming_entry_bit_concat14 = {FIRFilterStreaming_entry_bit_select13[28:0], FIRFilterStreaming_entry_bit_concat14_bit_select_operand_2[2:0]};
end
always @(*) begin
		FIRFilterStreaming_entry_sr_add17 = (FIRFilterStreaming_entry_11 + FIRFilterStreaming_entry_bit_concat16);
end
always @(*) begin
		FIRFilterStreaming_entry_sr_add18 = (FIRFilterStreaming_entry_bit_concat14 + FIRFilterStreaming_entry_sr_add17);
end
always @(*) begin
		FIRFilterStreaming_entry_bit_concat12 = {FIRFilterStreaming_entry_bit_select11[29:0], FIRFilterStreaming_entry_bit_concat12_bit_select_operand_2[1:0]};
end
always @(*) begin
		FIRFilterStreaming_entry_bit_concat10 = {FIRFilterStreaming_entry_bit_select9[28:0], FIRFilterStreaming_entry_bit_concat10_bit_select_operand_2[2:0]};
end
always @(*) begin
		FIRFilterStreaming_entry_sr_add21 = (FIRFilterStreaming_entry_bit_concat12 + FIRFilterStreaming_entry_bit_concat10);
end
always @(*) begin
		FIRFilterStreaming_entry_newEarly_newEarly_add_12 = (FIRFilterStreaming_entry_newEarly_newEarly_add_8_reg_stage1 + FIRFilterStreaming_entry_sr_add21_reg_stage1);
end
always @(*) begin
		FIRFilterStreaming_entry_bit_concat8 = {FIRFilterStreaming_entry_bit_select7[29:0], FIRFilterStreaming_entry_bit_concat8_bit_select_operand_2[1:0]};
end
always @(*) begin
		FIRFilterStreaming_entry_bit_concat6 = {FIRFilterStreaming_entry_bit_select5[28:0], FIRFilterStreaming_entry_bit_concat6_bit_select_operand_2[2:0]};
end
always @(*) begin
		FIRFilterStreaming_entry_sr_add24 = (FIRFilterStreaming_entry_13 + FIRFilterStreaming_entry_bit_concat8);
end
always @(*) begin
		FIRFilterStreaming_entry_sr_add25 = (FIRFilterStreaming_entry_bit_concat6 + FIRFilterStreaming_entry_sr_add24);
end
always @(*) begin
		FIRFilterStreaming_entry_newEarly_newEarly_add_13 = (FIRFilterStreaming_entry_sr_add18_reg_stage1 + FIRFilterStreaming_entry_sr_add25_reg_stage1);
end
always @(*) begin
		FIRFilterStreaming_entry_sr_negate24 = (32'd0 - FIRFilterStreaming_entry_14);
end
always @(*) begin
		FIRFilterStreaming_entry_bit_select3 = FIRFilterStreaming_entry_sr_negate24[30:0];
end
always @(*) begin
		FIRFilterStreaming_entry_bit_concat4 = {FIRFilterStreaming_entry_bit_select3[30:0], FIRFilterStreaming_entry_bit_concat4_bit_select_operand_2};
end
always @(*) begin
		FIRFilterStreaming_entry_bit_concat2 = {FIRFilterStreaming_entry_bit_select1[27:0], FIRFilterStreaming_entry_bit_concat2_bit_select_operand_2[3:0]};
end
always @(*) begin
		FIRFilterStreaming_entry_sr_add27 = (FIRFilterStreaming_entry_bit_concat4 + FIRFilterStreaming_entry_bit_concat2);
end
always @(*) begin
		FIRFilterStreaming_entry_newEarly_newEarly_newEarl = (FIRFilterStreaming_entry_sr_add13_reg_stage1 + FIRFilterStreaming_entry_sr_add27_reg_stage1);
end
always @(*) begin
		FIRFilterStreaming_entry_newCurOp_newEarly_newEarl = (FIRFilterStreaming_entry_newEarly_add_4_reg_stage1 + FIRFilterStreaming_entry_newEarly_newEarly_newEarl);
end
always @(*) begin
		FIRFilterStreaming_entry_newCurOp_newEarly_add_14 = (FIRFilterStreaming_entry_newCurOp_newEarly_newEarl_reg_stage2 + FIRFilterStreaming_entry_newEarly_newEarly_add_12_reg_stage2);
end
always @(*) begin
		FIRFilterStreaming_entry_sr_negate26 = (32'd0 - FIRFilterStreaming_entry_15);
end
always @(*) begin
		FIRFilterStreaming_entry_bit_concat = {FIRFilterStreaming_entry_bit_select[27:0], FIRFilterStreaming_entry_bit_concat_bit_select_operand_2[3:0]};
end
always @(*) begin
		FIRFilterStreaming_entry_sr_add28 = (FIRFilterStreaming_entry_sr_negate26 + FIRFilterStreaming_entry_bit_concat);
end
always @(*) begin
		FIRFilterStreaming_entry_newEarly_newEarly_newEarl_var0 = (FIRFilterStreaming_entry_newEarly_add_5_reg_stage1 + FIRFilterStreaming_entry_sr_add28_reg_stage1);
end
always @(*) begin
		FIRFilterStreaming_entry_newCurOp_newEarly_newEarl_var1 = (FIRFilterStreaming_entry_newEarly_newEarly_newEarl_var0 + FIRFilterStreaming_entry_newEarly_newEarly_add_9);
end
always @(*) begin
		FIRFilterStreaming_entry_newCurOp_newEarly_add_15 = (FIRFilterStreaming_entry_newCurOp_newEarly_newEarl_var1_reg_stage2 + FIRFilterStreaming_entry_newEarly_newEarly_add_13_reg_stage2);
end
always @(*) begin
		FIRFilterStreaming_entry_newCurOp_add_15 = (FIRFilterStreaming_entry_newCurOp_newEarly_add_14 + FIRFilterStreaming_entry_newCurOp_newEarly_add_15);
end
always @(*) begin
		FIRFilterStreaming_entry_cmp13 = (FIRFilterStreaming_entry_0 == 32'd0);
end
always @(*) begin
		FIRFilterStreaming_entry_cond = (FIRFilterStreaming_entry_cmp13_reg_stage3 ? 32'd0 : FIRFilterStreaming_entry_newCurOp_add_15_reg_stage3);
end
always @(posedge clk) begin
	if (reset) begin
		FIRFilterStreaming_previous_0_inferred_reg <= 32'd0;
	end
	if (FIRFilterStreaming_state_enable_0) begin
		FIRFilterStreaming_previous_0_inferred_reg <= FIRFilterStreaming_entry_15;
	end
end
always @(posedge clk) begin
	if (reset) begin
		FIRFilterStreaming_previous_1_inferred_reg <= 32'd0;
	end
	if (FIRFilterStreaming_state_enable_0) begin
		FIRFilterStreaming_previous_1_inferred_reg <= FIRFilterStreaming_entry_14;
	end
end
always @(posedge clk) begin
	if (reset) begin
		FIRFilterStreaming_previous_2_inferred_reg <= 32'd0;
	end
	if (FIRFilterStreaming_state_enable_0) begin
		FIRFilterStreaming_previous_2_inferred_reg <= FIRFilterStreaming_entry_13;
	end
end
always @(posedge clk) begin
	if (reset) begin
		FIRFilterStreaming_previous_3_inferred_reg <= 32'd0;
	end
	if (FIRFilterStreaming_state_enable_0) begin
		FIRFilterStreaming_previous_3_inferred_reg <= FIRFilterStreaming_entry_12;
	end
end
always @(posedge clk) begin
	if (reset) begin
		FIRFilterStreaming_previous_4_inferred_reg <= 32'd0;
	end
	if (FIRFilterStreaming_state_enable_0) begin
		FIRFilterStreaming_previous_4_inferred_reg <= FIRFilterStreaming_entry_11;
	end
end
always @(posedge clk) begin
	if (reset) begin
		FIRFilterStreaming_previous_5_inferred_reg <= 32'd0;
	end
	if (FIRFilterStreaming_state_enable_0) begin
		FIRFilterStreaming_previous_5_inferred_reg <= FIRFilterStreaming_entry_10;
	end
end
always @(posedge clk) begin
	if (reset) begin
		FIRFilterStreaming_previous_6_inferred_reg <= 32'd0;
	end
	if (FIRFilterStreaming_state_enable_0) begin
		FIRFilterStreaming_previous_6_inferred_reg <= FIRFilterStreaming_entry_9;
	end
end
always @(posedge clk) begin
	if (reset) begin
		FIRFilterStreaming_previous_7_inferred_reg <= 32'd0;
	end
	if (FIRFilterStreaming_state_enable_0) begin
		FIRFilterStreaming_previous_7_inferred_reg <= FIRFilterStreaming_entry_8;
	end
end
always @(posedge clk) begin
	if (reset) begin
		FIRFilterStreaming_previous_8_inferred_reg <= 32'd0;
	end
	if (FIRFilterStreaming_state_enable_0) begin
		FIRFilterStreaming_previous_8_inferred_reg <= FIRFilterStreaming_entry_7;
	end
end
always @(posedge clk) begin
	if (reset) begin
		FIRFilterStreaming_previous_9_inferred_reg <= 32'd0;
	end
	if (FIRFilterStreaming_state_enable_0) begin
		FIRFilterStreaming_previous_9_inferred_reg <= FIRFilterStreaming_entry_6;
	end
end
always @(posedge clk) begin
	if (reset) begin
		FIRFilterStreaming_previous_10_inferred_reg <= 32'd0;
	end
	if (FIRFilterStreaming_state_enable_0) begin
		FIRFilterStreaming_previous_10_inferred_reg <= FIRFilterStreaming_entry_5;
	end
end
always @(posedge clk) begin
	if (reset) begin
		FIRFilterStreaming_previous_11_inferred_reg <= 32'd0;
	end
	if (FIRFilterStreaming_state_enable_0) begin
		FIRFilterStreaming_previous_11_inferred_reg <= FIRFilterStreaming_entry_4;
	end
end
always @(posedge clk) begin
	if (reset) begin
		FIRFilterStreaming_previous_12_inferred_reg <= 32'd0;
	end
	if (FIRFilterStreaming_state_enable_0) begin
		FIRFilterStreaming_previous_12_inferred_reg <= FIRFilterStreaming_entry_3;
	end
end
always @(posedge clk) begin
	if (reset) begin
		FIRFilterStreaming_previous_13_inferred_reg <= 32'd0;
	end
	if (FIRFilterStreaming_state_enable_0) begin
		FIRFilterStreaming_previous_13_inferred_reg <= FIRFilterStreaming_entry_2;
	end
end
always @(posedge clk) begin
	if (reset) begin
		FIRFilterStreaming_previous_14_inferred_reg <= 32'd0;
	end
	if (FIRFilterStreaming_state_enable_0) begin
		FIRFilterStreaming_previous_14_inferred_reg <= FIRFilterStreaming_entry_1;
	end
end
always @(posedge clk) begin
	if (~(FIRFilterStreaming_state_stall_0)) begin
		FIRFilterStreaming_valid_bit_0 <= (FIRFilterStreaming_II_counter & start);
	end
	if (reset) begin
		FIRFilterStreaming_valid_bit_0 <= 1'd0;
	end
end
always @(*) begin
	FIRFilterStreaming_state_stall_0 = 1'd0;
	if (FIRFilterStreaming_state_stall_1) begin
		FIRFilterStreaming_state_stall_0 = 1'd1;
	end
	if ((FIRFilterStreaming_valid_bit_0 & ~(input_fifo_consumed_valid))) begin
		FIRFilterStreaming_state_stall_0 = 1'd1;
	end
end
always @(*) begin
	FIRFilterStreaming_state_enable_0 = (FIRFilterStreaming_valid_bit_0 & ~(FIRFilterStreaming_state_stall_0));
end
always @(posedge clk) begin
	if (~(FIRFilterStreaming_state_stall_1)) begin
		FIRFilterStreaming_valid_bit_1 <= FIRFilterStreaming_state_enable_0;
	end
	if (reset) begin
		FIRFilterStreaming_valid_bit_1 <= 1'd0;
	end
end
always @(*) begin
	FIRFilterStreaming_state_stall_1 = 1'd0;
	if (FIRFilterStreaming_state_stall_2) begin
		FIRFilterStreaming_state_stall_1 = 1'd1;
	end
end
always @(*) begin
	FIRFilterStreaming_state_enable_1 = (FIRFilterStreaming_valid_bit_1 & ~(FIRFilterStreaming_state_stall_1));
end
always @(posedge clk) begin
	if (~(FIRFilterStreaming_state_stall_2)) begin
		FIRFilterStreaming_valid_bit_2 <= FIRFilterStreaming_state_enable_1;
	end
	if (reset) begin
		FIRFilterStreaming_valid_bit_2 <= 1'd0;
	end
end
always @(*) begin
	FIRFilterStreaming_state_stall_2 = 1'd0;
	if (FIRFilterStreaming_state_stall_3) begin
		FIRFilterStreaming_state_stall_2 = 1'd1;
	end
end
always @(*) begin
	FIRFilterStreaming_state_enable_2 = (FIRFilterStreaming_valid_bit_2 & ~(FIRFilterStreaming_state_stall_2));
end
always @(posedge clk) begin
	if (~(FIRFilterStreaming_state_stall_3)) begin
		FIRFilterStreaming_valid_bit_3 <= FIRFilterStreaming_state_enable_2;
	end
	if (reset) begin
		FIRFilterStreaming_valid_bit_3 <= 1'd0;
	end
end
always @(*) begin
	FIRFilterStreaming_state_stall_3 = 1'd0;
	if ((((FIRFilterStreaming_valid_bit_3 & output_fifo_valid_to_sink) & ~(output_fifo_ready_from_sink)) & (output_fifo_FIRFilterStreaming_state_3_not_accessed_due_to_stall_a | output_fifo_FIRFilterStreaming_state_3_stalln_reg))) begin
		FIRFilterStreaming_state_stall_3 = 1'd1;
	end
end
always @(*) begin
	FIRFilterStreaming_state_enable_3 = (FIRFilterStreaming_valid_bit_3 & ~(FIRFilterStreaming_state_stall_3));
end
always @(posedge clk) begin
	FIRFilterStreaming_II_counter <= 1'd1;
end
always @(posedge clk) begin
	if (FIRFilterStreaming_state_enable_0) begin
		FIRFilterStreaming_entry_newEarly_add_4_reg_stage1 <= FIRFilterStreaming_entry_newEarly_add_4;
	end
end
always @(posedge clk) begin
	if (FIRFilterStreaming_state_enable_0) begin
		FIRFilterStreaming_entry_newEarly_add_5_reg_stage1 <= FIRFilterStreaming_entry_newEarly_add_5;
	end
end
always @(posedge clk) begin
	if (FIRFilterStreaming_state_enable_0) begin
		FIRFilterStreaming_entry_sr_add8_reg_stage1 <= FIRFilterStreaming_entry_sr_add8;
	end
end
always @(posedge clk) begin
	if (FIRFilterStreaming_state_enable_0) begin
		FIRFilterStreaming_entry_newEarly_newEarly_add_8_reg_stage1 <= FIRFilterStreaming_entry_newEarly_newEarly_add_8;
	end
end
always @(posedge clk) begin
	if (FIRFilterStreaming_state_enable_0) begin
		FIRFilterStreaming_entry_sr_add10_reg_stage1 <= FIRFilterStreaming_entry_sr_add10;
	end
end
always @(posedge clk) begin
	if (FIRFilterStreaming_state_enable_0) begin
		FIRFilterStreaming_entry_sr_add13_reg_stage1 <= FIRFilterStreaming_entry_sr_add13;
	end
end
always @(posedge clk) begin
	if (FIRFilterStreaming_state_enable_0) begin
		FIRFilterStreaming_entry_sr_add18_reg_stage1 <= FIRFilterStreaming_entry_sr_add18;
	end
end
always @(posedge clk) begin
	if (FIRFilterStreaming_state_enable_0) begin
		FIRFilterStreaming_entry_sr_add21_reg_stage1 <= FIRFilterStreaming_entry_sr_add21;
	end
end
always @(posedge clk) begin
	if (FIRFilterStreaming_state_enable_1) begin
		FIRFilterStreaming_entry_newEarly_newEarly_add_12_reg_stage2 <= FIRFilterStreaming_entry_newEarly_newEarly_add_12;
	end
end
always @(posedge clk) begin
	if (FIRFilterStreaming_state_enable_0) begin
		FIRFilterStreaming_entry_sr_add25_reg_stage1 <= FIRFilterStreaming_entry_sr_add25;
	end
end
always @(posedge clk) begin
	if (FIRFilterStreaming_state_enable_1) begin
		FIRFilterStreaming_entry_newEarly_newEarly_add_13_reg_stage2 <= FIRFilterStreaming_entry_newEarly_newEarly_add_13;
	end
end
always @(posedge clk) begin
	if (FIRFilterStreaming_state_enable_0) begin
		FIRFilterStreaming_entry_sr_add27_reg_stage1 <= FIRFilterStreaming_entry_sr_add27;
	end
end
always @(posedge clk) begin
	if (FIRFilterStreaming_state_enable_1) begin
		FIRFilterStreaming_entry_newCurOp_newEarly_newEarl_reg_stage2 <= FIRFilterStreaming_entry_newCurOp_newEarly_newEarl;
	end
end
always @(posedge clk) begin
	if (FIRFilterStreaming_state_enable_0) begin
		FIRFilterStreaming_entry_sr_add28_reg_stage1 <= FIRFilterStreaming_entry_sr_add28;
	end
end
always @(posedge clk) begin
	if (FIRFilterStreaming_state_enable_1) begin
		FIRFilterStreaming_entry_newCurOp_newEarly_newEarl_var1_reg_stage2 <= FIRFilterStreaming_entry_newCurOp_newEarly_newEarl_var1;
	end
end
always @(posedge clk) begin
	if (FIRFilterStreaming_state_enable_2) begin
		FIRFilterStreaming_entry_newCurOp_add_15_reg_stage3 <= FIRFilterStreaming_entry_newCurOp_add_15;
	end
end
always @(posedge clk) begin
	if (FIRFilterStreaming_state_enable_0) begin
		FIRFilterStreaming_entry_cmp13_reg_stage1 <= FIRFilterStreaming_entry_cmp13;
	end
end
always @(posedge clk) begin
	if (FIRFilterStreaming_state_enable_1) begin
		FIRFilterStreaming_entry_cmp13_reg_stage2 <= FIRFilterStreaming_entry_cmp13_reg_stage1;
	end
end
always @(posedge clk) begin
	if (FIRFilterStreaming_state_enable_2) begin
		FIRFilterStreaming_entry_cmp13_reg_stage3 <= FIRFilterStreaming_entry_cmp13_reg_stage2;
	end
end
always @(posedge clk) begin
	if (input_fifo_consumed_taken) begin
		input_fifo_consumed_valid <= 1'd0;
	end
	if ((input_fifo_ready_to_source & input_fifo_valid_from_source)) begin
		input_fifo_consumed_valid <= 1'd1;
	end
	if (reset) begin
		input_fifo_consumed_valid <= 1'd0;
	end
end
always @(posedge clk) begin
	if ((input_fifo_ready_to_source & input_fifo_valid_from_source)) begin
		input_fifo_consumed_data <= input_fifo_data_from_source;
	end
	if (reset) begin
		input_fifo_consumed_data <= 1'd0;
	end
end
always @(*) begin
	input_fifo_consumed_taken = 1'd0;
	if (FIRFilterStreaming_valid_bit_0) begin
		input_fifo_consumed_taken = ~(FIRFilterStreaming_state_stall_0);
	end
end
assign FIRFilterStreaming_entry_bit_concat38_bit_select_operand_2 = 1'd0;
assign FIRFilterStreaming_entry_bit_concat36_bit_select_operand_2 = 1'd0;
assign FIRFilterStreaming_entry_bit_concat34_bit_select_operand_2 = 2'd0;
assign FIRFilterStreaming_entry_bit_concat32_bit_select_operand_2 = 2'd0;
assign FIRFilterStreaming_entry_bit_concat30_bit_select_operand_2 = 1'd0;
assign FIRFilterStreaming_entry_bit_concat28_bit_select_operand_2 = 2'd0;
assign FIRFilterStreaming_entry_bit_concat26_bit_select_operand_2 = 3'd0;
assign FIRFilterStreaming_entry_bit_concat24_bit_select_operand_2 = 3'd0;
assign FIRFilterStreaming_entry_bit_concat22_bit_select_operand_2 = 3'd0;
assign FIRFilterStreaming_entry_bit_concat20_bit_select_operand_2 = 1'd0;
assign FIRFilterStreaming_entry_bit_concat18_bit_select_operand_2 = 3'd0;
assign FIRFilterStreaming_entry_bit_concat16_bit_select_operand_2 = 1'd0;
assign FIRFilterStreaming_entry_bit_concat14_bit_select_operand_2 = 3'd0;
assign FIRFilterStreaming_entry_bit_concat12_bit_select_operand_2 = 2'd0;
assign FIRFilterStreaming_entry_bit_concat10_bit_select_operand_2 = 3'd0;
assign FIRFilterStreaming_entry_bit_concat8_bit_select_operand_2 = 2'd0;
assign FIRFilterStreaming_entry_bit_concat6_bit_select_operand_2 = 3'd0;
assign FIRFilterStreaming_entry_bit_concat4_bit_select_operand_2 = 1'd0;
assign FIRFilterStreaming_entry_bit_concat2_bit_select_operand_2 = 4'd0;
assign FIRFilterStreaming_entry_bit_concat_bit_select_operand_2 = 4'd0;
always @(posedge clk) begin
	output_fifo_FIRFilterStreaming_state_3_not_accessed_due_to_stall_a <= ((FIRFilterStreaming_state_stall_3 & output_fifo_valid_to_sink) & ~(output_fifo_ready_from_sink));
end
always @(posedge clk) begin
	output_fifo_FIRFilterStreaming_state_3_stalln_reg <= ~(FIRFilterStreaming_state_stall_3);
end
always @(*) begin
	output_fifo_FIRFilterStreaming_state_3_enable_cond_a = (FIRFilterStreaming_valid_bit_3 & (output_fifo_FIRFilterStreaming_state_3_not_accessed_due_to_stall_a | output_fifo_FIRFilterStreaming_state_3_stalln_reg));
end
always @(posedge clk) begin
	finish <= FIRFilterStreaming_state_enable_3;
end
always @(*) begin
	input_fifo_ready_to_source = (~(input_fifo_consumed_valid) | input_fifo_consumed_taken);
	if (reset) begin
		input_fifo_ready_to_source = 1'd0;
	end
end
always @(*) begin
		output_fifo_data_to_sink = FIRFilterStreaming_entry_cond;
end
always @(*) begin
	output_fifo_valid_to_sink = 1'd0;
	if (output_fifo_FIRFilterStreaming_state_3_enable_cond_a) begin
		output_fifo_valid_to_sink = 1'd1;
	end
end

endmodule
